module mod_1 (
  input logic [2:0] in,
  output logic [2:0] out
);

assign out = in;
endmodule   // mod_1

