module mod1 (
  input logic  in,
  output logic  test
);

assign test = in;
endmodule   // mod1

