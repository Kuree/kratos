module module1(a, b, c, f);
output f;
input a, b, c;
// Description goes here
endmodule

// alternatively
module module2(input a, b, c, output f);
// Description goes here
endmodule