module mod (
  input logic [15:0] a [15:0],
  input logic [15:0] c,
  output logic b
);

endmodule   // mod
