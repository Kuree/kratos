module mod (
  input logic [15:0] a [15:0],
  output logic b,
  input logic [15:0] c
);

endmodule   // mod
