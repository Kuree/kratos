module mod (
  input logic [5:0] [3:0] in,
  output logic [5:0] [3:0] out
);

assign out = in;
endmodule   // mod

