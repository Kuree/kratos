module child(a, f);
input a;
output f;
endmodule
