module top (
  input logic  in,
  output logic  out
);

assign out = in;
endmodule   // top

