module mod (
  input logic [255:0] a,
  output logic b,
  input logic [15:0] c
);

endmodule   // mod
