`ifndef KRATOS_PACKED_STRUCT_PKG
`define KRATOS_PACKED_STRUCT_PKG
package packed_struct_pkg;
typedef struct packed {
    logic [15:0] read;
    logic [15:0] data;
} config_data;

endpackage
`endif
